module Register_File(clk,rst,Write_Enable,WD3,A1,A2,A3,RD1,RD2);
    input clk,rst,Write_Enable;
    input [4:0]A1,A2,A3;
    input [31:0]WD3;
    output [31:0]RD1,RD2;

    reg [31:0] Register [31:0];

    always @ (posedge clk)
    begin
        if(Write_Enable && (A3 != 5'd0))
            Register[A3] <= WD3;
    end

    assign RD1 = (~rst) ? 32'd0 : Register[A1];
    assign RD2 = (~rst) ? 32'd0 : Register[A2];

    
    integer i;
    initial begin
        for (i = 0; i < 32; i = i + 1)
            Register[i] = 32'b0;
    end

endmodule
